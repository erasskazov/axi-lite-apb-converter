`define AW_AXI  32 //axilite  address width
`define DW_AXI  32 //axilite  data    width  
`define AU_AXI  0  //axilite  user signals width
`define AW_APB  32 //apb4     address width                   
`define DW_APB  32 //apb4     data    width     
